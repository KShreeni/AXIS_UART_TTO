/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_top_axis_uart (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
//  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
    assign uio_out[7:3] = 0;
  assign uio_oe  = 8'b00000011;
    top_axis_uart #(.DATA_BITS(8)) dut(.clk(clk),.rst(rst_n),.axis_data(ui_in),.axis_valid(uio_in[2]),.axis_last(uio_in[3]),.m_axis_ready(uio_out[2]),.uart_tx(uio_out[0]),.rx_valid(uio_out[1]),.rx_data(uo_out));
  // List all unused inputs to prevent warnings
    wire _unused = &{ena, clk, rst_n, uio_in[7:4], uio_in[1:0], 1'b0};

endmodule
